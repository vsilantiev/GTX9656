------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.7
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : jesd204b_rx4_init.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module jesd204b_rx4_init
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity jesd204b_rx4_init is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";          -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;               -- Set to 1 for simulation
    STABLE_CLOCK_PERIOD                     : integer   := 10;               --Period of the stable clock driving this state-machine, unit is [ns]
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0                -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;

    --_________________________________________________________________________
    --GT0  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT0_DRPCLK_IN                           : in   std_logic;
    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT0_DRPEN_IN                            : in   std_logic;
    GT0_DRPRDY_OUT                          : out  std_logic;
    GT0_DRPWE_IN                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT0_GTPRXN_IN                           : in   std_logic;
    GT0_GTPRXP_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT0_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT0_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    GT0_RXLPMHFHOLD_IN                      : in   std_logic;
    GT0_RXLPMLFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT0_GTTXRESET_IN                        : in   std_logic;

    --GT1  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    GT1_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT1_DRPCLK_IN                           : in   std_logic;
    GT1_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT1_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT1_DRPEN_IN                            : in   std_logic;
    GT1_DRPRDY_OUT                          : out  std_logic;
    GT1_DRPWE_IN                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    GT1_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT1_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT1_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT1_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT1_RXUSRCLK_IN                         : in   std_logic;
    GT1_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT1_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT1_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT1_GTPRXN_IN                           : in   std_logic;
    GT1_GTPRXP_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT1_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT1_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    GT1_RXLPMHFHOLD_IN                      : in   std_logic;
    GT1_RXLPMLFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT1_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT1_GTRXRESET_IN                        : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT1_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT1_GTTXRESET_IN                        : in   std_logic;

    --GT2  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    GT2_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT2_DRPCLK_IN                           : in   std_logic;
    GT2_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT2_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT2_DRPEN_IN                            : in   std_logic;
    GT2_DRPRDY_OUT                          : out  std_logic;
    GT2_DRPWE_IN                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    GT2_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT2_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT2_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT2_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT2_RXUSRCLK_IN                         : in   std_logic;
    GT2_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT2_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT2_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT2_GTPRXN_IN                           : in   std_logic;
    GT2_GTPRXP_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT2_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT2_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    GT2_RXLPMHFHOLD_IN                      : in   std_logic;
    GT2_RXLPMLFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT2_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT2_GTRXRESET_IN                        : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT2_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT2_GTTXRESET_IN                        : in   std_logic;


    --____________________________COMMON PORTS________________________________
    ----------------- Common Block - GTPE2_COMMON Clocking Ports ---------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    -------------------------- Common Block - PLL Ports ------------------------
    GT0_PLL0LOCK_OUT                        : out  std_logic;
    GT0_PLL0LOCKDETCLK_IN                   : in   std_logic;
    GT0_PLL0RESET_IN                        : in   std_logic


);

end jesd204b_rx4_init;
    
architecture RTL of jesd204b_rx4_init is

--**************************Component Declarations*****************************


component jesd204b_rx4 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP    : string    := "FALSE" -- Set to 1 to speed up sim reset

);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
    GT0_DRP_BUSY_OUT                        : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT0_DRPCLK_IN                           : in   std_logic;
    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT0_DRPEN_IN                            : in   std_logic;
    GT0_DRPRDY_OUT                          : out  std_logic;
    GT0_DRPWE_IN                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT0_GTPRXN_IN                           : in   std_logic;
    GT0_GTPRXP_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT0_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT0_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    GT0_RXLPMHFHOLD_IN                      : in   std_logic;
    GT0_RXLPMLFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT0_TXPCSRESET_IN                       : in   std_logic;
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
    GT1_DRP_BUSY_OUT                        : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT1_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT1_DRPCLK_IN                           : in   std_logic;
    GT1_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT1_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT1_DRPEN_IN                            : in   std_logic;
    GT1_DRPRDY_OUT                          : out  std_logic;
    GT1_DRPWE_IN                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    GT1_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT1_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT1_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT1_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT1_RXUSRCLK_IN                         : in   std_logic;
    GT1_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT1_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT1_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT1_GTPRXN_IN                           : in   std_logic;
    GT1_GTPRXP_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT1_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT1_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    GT1_RXLPMHFHOLD_IN                      : in   std_logic;
    GT1_RXLPMLFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT1_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT1_GTRXRESET_IN                        : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT1_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT1_GTTXRESET_IN                        : in   std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT1_TXPCSRESET_IN                       : in   std_logic;
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
    GT2_DRP_BUSY_OUT                        : out  std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT2_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT2_DRPCLK_IN                           : in   std_logic;
    GT2_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT2_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT2_DRPEN_IN                            : in   std_logic;
    GT2_DRPRDY_OUT                          : out  std_logic;
    GT2_DRPWE_IN                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    GT2_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT2_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT2_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT2_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    GT2_RXUSRCLK_IN                         : in   std_logic;
    GT2_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT2_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT2_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT2_GTPRXN_IN                           : in   std_logic;
    GT2_GTPRXP_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT2_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT2_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    GT2_RXLPMHFHOLD_IN                      : in   std_logic;
    GT2_RXLPMLFHOLD_IN                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT2_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT2_GTRXRESET_IN                        : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT2_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT2_GTTXRESET_IN                        : in   std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT2_TXPCSRESET_IN                       : in   std_logic;
   

    --____________________________COMMON PORTS________________________________
    ----------------- Common Block - GTPE2_COMMON Clocking Ports ---------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    -------------------------- Common Block - PLL Ports ------------------------
    GT0_PLL0LOCK_OUT                        : out  std_logic;
    GT0_PLL0LOCKDETCLK_IN                   : in   std_logic;
    GT0_PLL0REFCLKLOST_OUT                  : out  std_logic;
    GT0_PLL0RESET_IN                        : in   std_logic


);
end component;

component jesd204b_rx4_TX_STARTUP_FSM
  Generic(
           GT_TYPE                  : string := "GTX";
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
            TX_PLL0_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_PLL0_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient              
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           TXUSERCLK                : in  STD_LOGIC;              --TXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;              --User Reset, can be pulled any time
           PLL0REFCLKLOST           : in  STD_LOGIC;              --PLL0 Reference-clock for the GT is lost
           PLL1REFCLKLOST           : in  STD_LOGIC;              --PLL1 Reference-clock for the GT is lost
           PLL0LOCK                 : in  STD_LOGIC;              --Lock Detect from the PLL0 of the GT
           PLL1LOCK                 : in  STD_LOGIC;              --Lock Detect from the PLL1 of the GT
           TXRESETDONE              : in  STD_LOGIC;      
           MMCM_LOCK                : in  STD_LOGIC;      
           GTTXRESET                : out STD_LOGIC:='0';      
           MMCM_RESET               : out STD_LOGIC:='0';      
           PLL0_RESET               : out STD_LOGIC:='0';        --Reset PLL0
           PLL1_RESET               : out STD_LOGIC:='0';        --Reset PLL1
           TX_FSM_RESET_DONE        : out STD_LOGIC:='0';        --Reset-sequence has sucessfully been finished.
           TXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC:='0';
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';
           PHALIGNMENT_DONE         : in  STD_LOGIC;
           
           RETRY_COUNTER            : out  STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;

component jesd204b_rx4_RX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           GT_TYPE                  : string := "GTX";
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_PLL0_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_PLL0_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient                         
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;        --Stable Clock, either a stable clock from the PCB
                                                            --or reference-clock present at startup.
           RXUSERCLK                : in  STD_LOGIC;        --RXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;        --User Reset, can be pulled any time
           PLL0REFCLKLOST           : in  STD_LOGIC;        --PLL0 Reference-clock for the GT is lost
           PLL1REFCLKLOST           : in  STD_LOGIC;        --PLL1 Reference-clock for the GT is lost
           PLL0LOCK                 : in  STD_LOGIC;        --Lock Detect from the PLL0 of the GT
           PLL1LOCK                 : in  STD_LOGIC;        --Lock Detect from the PLL1 of the GT
           RXRESETDONE              : in  STD_LOGIC;
           MMCM_LOCK                : in  STD_LOGIC;
           RECCLK_STABLE            : in  STD_LOGIC;
           RECCLK_MONITOR_RESTART   : in  STD_LOGIC;
           DATA_VALID               : in  STD_LOGIC;
           TXUSERRDY                : in  STD_LOGIC;       --TXUSERRDY from GT 
           DONT_RESET_ON_DATA_ERROR : in  STD_LOGIC;
           GTRXRESET                : out STD_LOGIC:='0';
           MMCM_RESET               : out STD_LOGIC:='0';
           PLL0_RESET               : out STD_LOGIC:='0';  --Reset PLL0 (only if RX uses PLL0)
           PLL1_RESET               : out STD_LOGIC:='0';  --Reset PLL1 (only if RX uses PLL1)
           RX_FSM_RESET_DONE        : out STD_LOGIC:='0';  --Reset-sequence has sucessfully been finished.
           RXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC;
           PHALIGNMENT_DONE         : in  STD_LOGIC; 
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';           
           RETRY_COUNTER            : out STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;






  function get_cdrlock_time(is_sim : in integer) return integer is
    variable lock_time: integer;
  begin
    if (is_sim = 1) then
      lock_time := 1000;
    else
      lock_time := 50000 / integer(3.072); --Typical CDR lock time is 50,000UI as per DS183
    end if;
    return lock_time;
  end function;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    constant RX_CDRLOCK_TIME      : integer := get_cdrlock_time(EXAMPLE_SIMULATION);       -- 200us
    constant WAIT_TIME_CDRLOCK    : integer := RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      -- 200 us time-out

    -------------------------- GT Wrapper Wires ------------------------------
    signal   gt0_txresetdone_i               : std_logic;
    signal   gt0_rxresetdone_i               : std_logic;
    signal   gt0_gttxreset_i                 : std_logic;
    signal   gt0_gttxreset_t                 : std_logic;
    signal   gt0_gtrxreset_i                 : std_logic;
    signal   gt0_gtrxreset_t                 : std_logic;
    signal   gt0_txpcsreset_i                : std_logic;
    signal   gt0_txuserrdy_i                 : std_logic;
    signal   gt0_txuserrdy_t                 : std_logic;
    signal   gt0_rxuserrdy_i                 : std_logic;
    signal   gt0_rxuserrdy_t                 : std_logic;



    signal   gt1_txresetdone_i               : std_logic;
    signal   gt1_rxresetdone_i               : std_logic;
    signal   gt1_gttxreset_i                 : std_logic;
    signal   gt1_gttxreset_t                 : std_logic;
    signal   gt1_gtrxreset_i                 : std_logic;
    signal   gt1_gtrxreset_t                 : std_logic;
    signal   gt1_txpcsreset_i                : std_logic;
    signal   gt1_txuserrdy_i                 : std_logic;
    signal   gt1_txuserrdy_t                 : std_logic;
    signal   gt1_rxuserrdy_i                 : std_logic;
    signal   gt1_rxuserrdy_t                 : std_logic;



    signal   gt2_txresetdone_i               : std_logic;
    signal   gt2_rxresetdone_i               : std_logic;
    signal   gt2_gttxreset_i                 : std_logic;
    signal   gt2_gttxreset_t                 : std_logic;
    signal   gt2_gtrxreset_i                 : std_logic;
    signal   gt2_gtrxreset_t                 : std_logic;
    signal   gt2_txpcsreset_i                : std_logic;
    signal   gt2_txuserrdy_i                 : std_logic;
    signal   gt2_txuserrdy_t                 : std_logic;
    signal   gt2_rxuserrdy_i                 : std_logic;
    signal   gt2_rxuserrdy_t                 : std_logic;




    signal   gt0_pll0reset_i                 : std_logic;
    signal   gt0_pll0reset_t                 : std_logic;
    signal   gt0_pll0refclklost_i            : std_logic;
    signal   gt0_pll0lock_i                  : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_vcc_i                   : std_logic;

    signal   gt0_rxoutclk_i                  : std_logic;
    signal   gt0_recclk_stable_i             : std_logic;

    signal   gt1_rxoutclk_i                  : std_logic;
    signal   gt1_recclk_stable_i             : std_logic;

    signal   gt2_rxoutclk_i                  : std_logic;
    signal   gt2_recclk_stable_i             : std_logic;






    signal   rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;
    signal      rx_cdrlocked                    : std_logic;


 


--**************************** Main Body of Code *******************************
begin
    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_vcc_i                                <= '1';

    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    jesd204b_rx4_i : jesd204b_rx4
    generic map
    (
        WRAPPER_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP
    )
    port map
    (
        GT0_DRP_BUSY_OUT                =>      open,
  
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X0Y1)

        ---------------------------- Channel - DRP Ports  --------------------------
        GT0_DRPADDR_IN                  =>      GT0_DRPADDR_IN,
        GT0_DRPCLK_IN                   =>      GT0_DRPCLK_IN,
        GT0_DRPDI_IN                    =>      GT0_DRPDI_IN,
        GT0_DRPDO_OUT                   =>      GT0_DRPDO_OUT,
        GT0_DRPEN_IN                    =>      GT0_DRPEN_IN,
        GT0_DRPRDY_OUT                  =>      GT0_DRPRDY_OUT,
        GT0_DRPWE_IN                    =>      GT0_DRPWE_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        GT0_RXUSERRDY_IN                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT0_EYESCANDATAERROR_OUT        =>      GT0_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT0_RXCDRLOCK_OUT               =>      GT0_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT0_RXDATA_OUT                  =>      GT0_RXDATA_OUT,
        GT0_RXUSRCLK_IN                 =>      GT0_RXUSRCLK_IN,
        GT0_RXUSRCLK2_IN                =>      GT0_RXUSRCLK2_IN,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT0_RXCHARISCOMMA_OUT           =>      GT0_RXCHARISCOMMA_OUT,
        GT0_RXCHARISK_OUT               =>      GT0_RXCHARISK_OUT,
        GT0_RXDISPERR_OUT               =>      GT0_RXDISPERR_OUT,
        GT0_RXNOTINTABLE_OUT            =>      GT0_RXNOTINTABLE_OUT,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT0_GTPRXN_IN                   =>      GT0_GTPRXN_IN,
        GT0_GTPRXP_IN                   =>      GT0_GTPRXP_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT0_RXMCOMMAALIGNEN_IN          =>      GT0_RXMCOMMAALIGNEN_IN,
        GT0_RXPCOMMAALIGNEN_IN          =>      GT0_RXPCOMMAALIGNEN_IN,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        GT0_RXLPMHFHOLD_IN              =>      GT0_RXLPMHFHOLD_IN,
        GT0_RXLPMLFHOLD_IN              =>      GT0_RXLPMLFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT0_RXOUTCLK_OUT                =>      gt0_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT0_GTRXRESET_IN                =>      gt0_gtrxreset_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT0_RXRESETDONE_OUT             =>      gt0_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT0_GTTXRESET_IN                =>      gt0_gttxreset_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT0_TXPCSRESET_IN               =>      gt0_txpcsreset_i,


        GT1_DRP_BUSY_OUT                =>      open,
  
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X0Y2)

        ---------------------------- Channel - DRP Ports  --------------------------
        GT1_DRPADDR_IN                  =>      GT1_DRPADDR_IN,
        GT1_DRPCLK_IN                   =>      GT1_DRPCLK_IN,
        GT1_DRPDI_IN                    =>      GT1_DRPDI_IN,
        GT1_DRPDO_OUT                   =>      GT1_DRPDO_OUT,
        GT1_DRPEN_IN                    =>      GT1_DRPEN_IN,
        GT1_DRPRDY_OUT                  =>      GT1_DRPRDY_OUT,
        GT1_DRPWE_IN                    =>      GT1_DRPWE_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        GT1_RXUSERRDY_IN                =>      gt1_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT1_EYESCANDATAERROR_OUT        =>      GT1_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT1_RXCDRLOCK_OUT               =>      GT1_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT1_RXDATA_OUT                  =>      GT1_RXDATA_OUT,
        GT1_RXUSRCLK_IN                 =>      GT1_RXUSRCLK_IN,
        GT1_RXUSRCLK2_IN                =>      GT1_RXUSRCLK2_IN,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT1_RXCHARISCOMMA_OUT           =>      GT1_RXCHARISCOMMA_OUT,
        GT1_RXCHARISK_OUT               =>      GT1_RXCHARISK_OUT,
        GT1_RXDISPERR_OUT               =>      GT1_RXDISPERR_OUT,
        GT1_RXNOTINTABLE_OUT            =>      GT1_RXNOTINTABLE_OUT,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT1_GTPRXN_IN                   =>      GT1_GTPRXN_IN,
        GT1_GTPRXP_IN                   =>      GT1_GTPRXP_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT1_RXMCOMMAALIGNEN_IN          =>      GT1_RXMCOMMAALIGNEN_IN,
        GT1_RXPCOMMAALIGNEN_IN          =>      GT1_RXPCOMMAALIGNEN_IN,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        GT1_RXLPMHFHOLD_IN              =>      GT1_RXLPMHFHOLD_IN,
        GT1_RXLPMLFHOLD_IN              =>      GT1_RXLPMLFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT1_RXOUTCLK_OUT                =>      gt1_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT1_GTRXRESET_IN                =>      gt1_gtrxreset_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT1_RXRESETDONE_OUT             =>      gt1_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT1_GTTXRESET_IN                =>      gt1_gttxreset_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT1_TXPCSRESET_IN               =>      gt1_txpcsreset_i,


        GT2_DRP_BUSY_OUT                =>      open,
  
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X0Y3)

        ---------------------------- Channel - DRP Ports  --------------------------
        GT2_DRPADDR_IN                  =>      GT2_DRPADDR_IN,
        GT2_DRPCLK_IN                   =>      GT2_DRPCLK_IN,
        GT2_DRPDI_IN                    =>      GT2_DRPDI_IN,
        GT2_DRPDO_OUT                   =>      GT2_DRPDO_OUT,
        GT2_DRPEN_IN                    =>      GT2_DRPEN_IN,
        GT2_DRPRDY_OUT                  =>      GT2_DRPRDY_OUT,
        GT2_DRPWE_IN                    =>      GT2_DRPWE_IN,
        --------------------- RX Initialization and Reset Ports --------------------
        GT2_RXUSERRDY_IN                =>      gt2_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT2_EYESCANDATAERROR_OUT        =>      GT2_EYESCANDATAERROR_OUT,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT2_RXCDRLOCK_OUT               =>      GT2_RXCDRLOCK_OUT,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT2_RXDATA_OUT                  =>      GT2_RXDATA_OUT,
        GT2_RXUSRCLK_IN                 =>      GT2_RXUSRCLK_IN,
        GT2_RXUSRCLK2_IN                =>      GT2_RXUSRCLK2_IN,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT2_RXCHARISCOMMA_OUT           =>      GT2_RXCHARISCOMMA_OUT,
        GT2_RXCHARISK_OUT               =>      GT2_RXCHARISK_OUT,
        GT2_RXDISPERR_OUT               =>      GT2_RXDISPERR_OUT,
        GT2_RXNOTINTABLE_OUT            =>      GT2_RXNOTINTABLE_OUT,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT2_GTPRXN_IN                   =>      GT2_GTPRXN_IN,
        GT2_GTPRXP_IN                   =>      GT2_GTPRXP_IN,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT2_RXMCOMMAALIGNEN_IN          =>      GT2_RXMCOMMAALIGNEN_IN,
        GT2_RXPCOMMAALIGNEN_IN          =>      GT2_RXPCOMMAALIGNEN_IN,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        GT2_RXLPMHFHOLD_IN              =>      GT2_RXLPMHFHOLD_IN,
        GT2_RXLPMLFHOLD_IN              =>      GT2_RXLPMLFHOLD_IN,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT2_RXOUTCLK_OUT                =>      gt2_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT2_GTRXRESET_IN                =>      gt2_gtrxreset_i,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT2_RXRESETDONE_OUT             =>      gt2_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT2_GTTXRESET_IN                =>      gt2_gttxreset_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT2_TXPCSRESET_IN               =>      gt2_txpcsreset_i,




    --____________________________COMMON PORTS________________________________
        ----------------- Common Block - GTPE2_COMMON Clocking Ports ---------------
        GT0_GTREFCLK0_IN                =>      GT0_GTREFCLK0_IN,
        -------------------------- Common Block - PLL Ports ------------------------
        GT0_PLL0LOCK_OUT                =>      gt0_pll0lock_i,
        GT0_PLL0LOCKDETCLK_IN           =>      GT0_PLL0LOCKDETCLK_IN,
        GT0_PLL0REFCLKLOST_OUT          =>      gt0_pll0refclklost_i,
        GT0_PLL0RESET_IN                =>      gt0_pll0reset_i

    );

    gt0_txpcsreset_i                             <= tied_to_ground_i;
    gt1_txpcsreset_i                             <= tied_to_ground_i;
    gt2_txpcsreset_i                             <= tied_to_ground_i;





    GT0_RXRESETDONE_OUT                          <= gt0_rxresetdone_i;
    GT0_RXOUTCLK_OUT                             <= gt0_rxoutclk_i;
    GT1_RXRESETDONE_OUT                          <= gt1_rxresetdone_i;
    GT1_RXOUTCLK_OUT                             <= gt1_rxoutclk_i;
    GT2_RXRESETDONE_OUT                          <= gt2_rxresetdone_i;
    GT2_RXOUTCLK_OUT                             <= gt2_rxoutclk_i;
    GT0_PLL0LOCK_OUT                             <= gt0_pll0lock_i;

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    gt0_gttxreset_i                              <= GT0_GTTXRESET_IN or gt0_gttxreset_t;
    gt0_gtrxreset_i                              <= GT0_GTRXRESET_IN or gt0_gtrxreset_t;
    gt0_rxuserrdy_i                              <= GT0_RXUSERRDY_IN or gt0_rxuserrdy_t;
    gt1_gttxreset_i                              <= GT1_GTTXRESET_IN or gt1_gttxreset_t;
    gt1_gtrxreset_i                              <= GT1_GTRXRESET_IN or gt1_gtrxreset_t;
    gt1_rxuserrdy_i                              <= GT1_RXUSERRDY_IN or gt1_rxuserrdy_t;
    gt2_gttxreset_i                              <= GT2_GTTXRESET_IN or gt2_gttxreset_t;
    gt2_gtrxreset_i                              <= GT2_GTRXRESET_IN or gt2_gtrxreset_t;
    gt2_rxuserrdy_i                              <= GT2_RXUSERRDY_IN or gt2_rxuserrdy_t;
    gt0_pll0reset_i                              <= GT0_PLL0RESET_IN or gt0_pll0reset_t;
end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate
    gt0_gttxreset_i                              <= gt0_gttxreset_t;
    gt0_gtrxreset_i                              <= gt0_gtrxreset_t;
    gt0_txuserrdy_i                              <= gt0_txuserrdy_t;
    gt0_rxuserrdy_i                              <= gt0_rxuserrdy_t;
    gt1_gttxreset_i                              <= gt1_gttxreset_t;
    gt1_gtrxreset_i                              <= gt1_gtrxreset_t;
    gt1_txuserrdy_i                              <= gt1_txuserrdy_t;
    gt1_rxuserrdy_i                              <= gt1_rxuserrdy_t;
    gt2_gttxreset_i                              <= gt2_gttxreset_t;
    gt2_gtrxreset_i                              <= gt2_gtrxreset_t;
    gt2_txuserrdy_i                              <= gt2_txuserrdy_t;
    gt2_rxuserrdy_i                              <= gt2_rxuserrdy_t;
    gt0_pll0reset_i                              <= gt0_pll0reset_t;
end generate no_chipscope;






gt0_rxresetfsm_i:  jesd204b_rx4_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTP", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_PLL0_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_PLL0_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT0_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        PLL0REFCLKLOST                  =>      gt0_pll0refclklost_i,
        PLL0LOCK                        =>      gt0_pll0lock_i,
        PLL1REFCLKLOST                  =>      tied_to_ground_i,
        PLL1LOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt0_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT0_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt0_gtrxreset_t,
        MMCM_RESET                      =>      open,
        PLL0_RESET                      =>      gt0_pll0reset_t,
        PLL1_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT0_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt0_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt1_rxresetfsm_i:  jesd204b_rx4_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTP", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_PLL0_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_PLL0_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT1_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        PLL0REFCLKLOST                  =>      gt0_pll0refclklost_i,
        PLL0LOCK                        =>      gt0_pll0lock_i,
        PLL1REFCLKLOST                  =>      tied_to_ground_i,
        PLL1LOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt1_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt1_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT1_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt1_gtrxreset_t,
        MMCM_RESET                      =>      open,
        PLL0_RESET                      =>      open,
        PLL1_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT1_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt1_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt2_rxresetfsm_i:  jesd204b_rx4_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           GT_TYPE                  => "GTP", --GTX or GTH or GTP
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_PLL0_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_PLL0_USED             => TRUE,                         -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT2_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        PLL0REFCLKLOST                  =>      gt0_pll0refclklost_i,
        PLL0LOCK                        =>      gt0_pll0lock_i,
        PLL1REFCLKLOST                  =>      tied_to_ground_i,
        PLL1LOCK                        =>      tied_to_vcc_i,
        RXRESETDONE                     =>      gt2_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt2_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT2_DATA_VALID_IN,
        TXUSERRDY                       =>      tied_to_vcc_i,
        GTRXRESET                       =>      gt2_gtrxreset_t,
        MMCM_RESET                      =>      open,
        PLL0_RESET                      =>      open,
        PLL1_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT2_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt2_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );



  cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt0_gtrxreset_i = '1') then
          rx_cdrlocked       <= '0';
          rx_cdrlock_counter <=  0                        after DLY;
        elsif (rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          rx_cdrlocked       <= '1';
          rx_cdrlock_counter <= rx_cdrlock_counter        after DLY;
        else
          rx_cdrlock_counter <= rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

gt0_recclk_stable_i                          <= rx_cdrlocked;
gt1_recclk_stable_i                          <= rx_cdrlocked;
gt2_recclk_stable_i                          <= rx_cdrlocked;







end RTL;


